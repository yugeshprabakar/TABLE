//module declaration
module ksa64x64(x,y,sum,cin,cout);
//port declaration
input[63:0]x,y;
output[63:0]sum;
input [31:0]cin;
output cout;
//internal wire
wire[63:0]g1,p1,g2;
wire[64:2]g3;
wire[64:8]p4;
wire[64:4]p3;
wire[63:1]p2;
wire[64:4]g4;
wire[64:8]g5;
wire[64:16]p5;
wire[64:16]g6;
wire[63:32]g7;
wire[64:32]p6;
//gate instantiation
//level1
gray_cell l0A(cin[0],p1[0],g1[0],g2[0]);
black_cell l1A(g1[0],p1[1],g1[1],p1[0],g2[1],p2[1]);
black_cell l2A(g1[1],p1[2],g1[2],p1[1],g2[2],p2[2]);
black_cell l3A(g1[2],p1[3],g1[3],p1[2],g2[3],p2[3]);
black_cell l4A(g1[3],p1[4],g1[4],p1[3],g2[4],p2[4]);
black_cell l5A(g1[4],p1[5],g1[5],p1[4],g2[5],p2[5]);
black_cell l6A(g1[5],p1[6],g1[6],p1[5],g2[6],p2[6]);
black_cell l7A(g1[6],p1[7],g1[7],p1[6],g2[7],p2[7]);
black_cell l8A(g1[7],p1[8],g1[8],p1[7],g2[8],p2[8]);
black_cell l9A(g1[8],p1[9],g1[9],p1[8],g2[9],p2[9]);
black_cell l10A(g1[9],p1[10],g1[10],p1[9],g2[10],p2[10]);
black_cell l11A(g1[10],p1[11],g1[11],p1[10],g2[11],p2[11]);
black_cell l12A(g1[11],p1[12],g1[12],p1[11],g2[12],p2[12]);
black_cell l13A(g1[12],p1[13],g1[13],p1[12],g2[13],p2[13]);
black_cell l14A(g1[13],p1[14],g1[14],p1[13],g2[14],p2[14]);
black_cell l15A(g1[14],p1[15],g1[15],p1[14],g2[15],p2[15]);
black_cell l16A(g1[15],p1[16],g1[16],p1[15],g2[16],p2[16]);
black_cell l17A(g1[16],p1[17],g1[17],p1[16],g2[17],p2[17]);
black_cell l18A(g1[17],p1[18],g1[18],p1[17],g2[18],p2[18]);
black_cell l19A(g1[18],p1[19],g1[19],p1[18],g2[19],p2[19]);
black_cell l20A(g1[19],p1[20],g1[20],p1[19],g2[20],p2[20]);
black_cell l21A(g1[20],p1[21],g1[21],p1[20],g2[21],p2[21]);
black_cell l22A(g1[21],p1[22],g1[22],p1[21],g2[22],p2[22]);
black_cell l23A(g1[22],p1[23],g1[23],p1[22],g2[23],p2[23]);
black_cell l24A(g1[23],p1[24],g1[24],p1[23],g2[24],p2[24]);
black_cell l25A(g1[24],p1[25],g1[25],p1[24],g2[25],p2[25]);
black_cell l26A(g1[25],p1[26],g1[26],p1[25],g2[26],p2[26]);
black_cell l27A(g1[26],p1[27],g1[27],p1[26],g2[27],p2[27]);
black_cell l28A(g1[27],p1[28],g1[28],p1[27],g2[28],p2[28]);
black_cell l29A(g1[28],p1[29],g1[29],p1[28],g2[29],p2[29]);
black_cell l30A(g1[29],p1[30],g1[30],p1[29],g2[30],p2[30]);
black_cell l31A(g1[30],p1[31],g1[31],p1[30],g2[31],p2[31]);
black_cell l32A(g1[31],p1[32],g1[32],p1[31],g2[32],p2[32]);
black_cell l33A(g1[32],p1[33],g1[33],p1[32],g2[33],p2[33]);
black_cell l34A(g1[33],p1[34],g1[34],p1[33],g2[34],p2[34]);
black_cell l35A(g1[34],p1[35],g1[35],p1[34],g2[35],p2[35]);
black_cell l36A(g1[35],p1[36],g1[36],p1[35],g2[36],p2[36]);
black_cell l37A(g1[36],p1[37],g1[37],p1[36],g2[37],p2[37]);
black_cell l38A(g1[37],p1[38],g1[38],p1[37],g2[38],p2[38]);
black_cell l39A(g1[38],p1[39],g1[39],p1[38],g2[39],p2[39]);
black_cell l40A(g1[39],p1[40],g1[40],p1[39],g2[40],p2[40]);
black_cell l41A(g1[40],p1[41],g1[41],p1[40],g2[41],p2[41]);
black_cell l42A(g1[41],p1[42],g1[42],p1[41],g2[42],p2[42]);
black_cell l43A(g1[42],p1[43],g1[43],p1[42],g2[43],p2[43]);
black_cell l44A(g1[43],p1[44],g1[44],p1[43],g2[44],p2[44]);
black_cell l45A(g1[44],p1[45],g1[45],p1[44],g2[45],p2[45]);
black_cell l46A(g1[45],p1[46],g1[46],p1[45],g2[46],p2[46]);
black_cell l47A(g1[46],p1[47],g1[47],p1[46],g2[47],p2[47]);
black_cell l48A(g1[47],p1[48],g1[48],p1[47],g2[48],p2[48]);
black_cell l49A(g1[48],p1[49],g1[49],p1[48],g2[49],p2[49]);
black_cell l50A(g1[49],p1[50],g1[50],p1[49],g2[50],p2[50]);
black_cell l51A(g1[50],p1[51],g1[51],p1[50],g2[51],p2[51]);
black_cell l52A(g1[51],p1[52],g1[52],p1[51],g2[52],p2[52]);
black_cell l53A(g1[52],p1[53],g1[53],p1[52],g2[53],p2[53]);
black_cell l54A(g1[53],p1[54],g1[54],p1[53],g2[54],p2[54]);
black_cell l55A(g1[54],p1[55],g1[55],p1[54],g2[55],p2[55]);
black_cell l56A(g1[55],p1[56],g1[56],p1[55],g2[56],p2[56]);
black_cell l57A(g1[56],p1[57],g1[57],p1[56],g2[57],p2[57]);
black_cell l58A(g1[57],p1[58],g1[58],p1[57],g2[58],p2[58]);
black_cell l59A(g1[58],p1[59],g1[59],p1[58],g2[59],p2[59]);
black_cell l60A(g1[59],p1[60],g1[60],p1[59],g2[60],p2[60]);
black_cell l61A(g1[60],p1[61],g1[61],p1[60],g2[61],p2[61]);
black_cell l62A(g1[61],p1[62],g1[62],p1[61],g2[62],p2[62]);
black_cell l63A(g1[62],p1[63],g1[63],p1[62],g2[63],p2[63]);
//level
gray_cell l1B(cin[0],p2[1],g2[1],g3[2]);
gray_cell l2B(g2[0],p2[2],g2[2],g3[3]);
black_cell l3B(g2[1],p2[3],g2[3],p2[1],g3[4],p3[4]);
black_cell l4B(g2[2],p2[4],g2[4],p2[2],g3[5],p3[5]);
black_cell l5B(g2[3],p2[5],g2[5],p2[3],g3[6],p3[6]);
black_cell l6B(g2[4],p2[6],g2[6],p2[4],g3[7],p3[7]);
black_cell l7B(g2[5],p2[7],g2[7],p2[5],g3[8],p3[8]);
black_cell l8B(g2[6],p2[8],g2[8],p2[6],g3[9],p3[9]);
black_cell l9B(g2[7],p2[9],g2[9],p2[7],g3[10],p3[10]);
black_cell l10B(g2[8],p2[10],g2[10],p2[8],g3[11],p3[11]);
black_cell l11B(g2[9],p2[11],g2[11],p2[9],g3[12],p3[12]);
black_cell l12B(g2[10],p2[12],g2[12],p2[10],g3[13],p3[13]);
black_cell l13B(g2[11],p2[13],g2[13],p2[11],g3[14],p3[14]);
black_cell l14B(g2[12],p2[14],g2[14],p2[12],g3[15],p3[15]);
black_cell l15B(g2[13],p2[15],g2[15],p2[13],g3[16],p3[16]);
black_cell l16B(g2[14],p2[16],g2[16],p2[14],g3[17],p3[17]);
black_cell l17B(g2[15],p2[17],g2[17],p2[15],g3[18],p3[18]);
black_cell l18B(g2[16],p2[18],g2[18],p2[16],g3[19],p3[19]);
black_cell l19B(g2[17],p2[19],g2[19],p2[17],g3[20],p3[20]);
black_cell l20B(g2[18],p2[20],g2[20],p2[18],g3[21],p3[21]);
black_cell l21B(g2[19],p2[21],g2[21],p2[19],g3[22],p3[22]);
black_cell l22B(g2[20],p2[22],g2[22],p2[20],g3[23],p3[23]);
black_cell l23B(g2[21],p2[23],g2[23],p2[21],g3[24],p3[24]);
black_cell l24B(g2[22],p2[24],g2[24],p2[22],g3[25],p3[25]);
black_cell l25B(g2[23],p2[25],g2[25],p2[23],g3[26],p3[26]);
black_cell l26B(g2[24],p2[26],g2[26],p2[24],g3[27],p3[27]);
black_cell l27B(g2[25],p2[27],g2[27],p2[25],g3[28],p3[28]);
black_cell l28B(g2[26],p2[28],g2[28],p2[26],g3[29],p3[29]);
black_cell l29B(g2[27],p2[29],g2[29],p2[27],g3[30],p3[30]);
black_cell l30B(g2[28],p2[30],g2[30],p2[28],g3[31],p3[31]);
black_cell l31B(g2[29],p2[31],g2[31],p2[29],g3[32],p3[32]);
black_cell l32B(g2[30],p2[32],g2[32],p2[30],g3[33],p3[33]);
black_cell l33B(g2[31],p2[33],g2[33],p2[31],g3[34],p3[34]);
black_cell l34B(g2[32],p2[34],g2[34],p2[32],g3[35],p3[35]);
black_cell l35B(g2[33],p2[35],g2[35],p2[33],g3[36],p3[36]);
black_cell l36B(g2[34],p2[36],g2[36],p2[34],g3[37],p3[37]);
black_cell l37B(g2[35],p2[37],g2[37],p2[35],g3[38],p3[38]);
black_cell l38B(g2[36],p2[38],g2[38],p2[36],g3[39],p3[39]);
black_cell l39B(g2[37],p2[39],g2[39],p2[37],g3[40],p3[40]);
black_cell l40B(g2[38],p2[40],g2[40],p2[38],g3[41],p3[41]);
black_cell l41B(g2[39],p2[41],g2[41],p2[39],g3[42],p3[42]);
black_cell l42B(g2[40],p2[42],g2[42],p2[40],g3[43],p3[43]);
black_cell l43B(g2[41],p2[43],g2[43],p2[41],g3[44],p3[44]);
black_cell l44B(g2[42],p2[44],g2[44],p2[42],g3[45],p3[45]);
black_cell l45B(g2[43],p2[45],g2[45],p2[43],g3[46],p3[46]);
black_cell l46B(g2[44],p2[46],g2[46],p2[44],g3[47],p3[47]);
black_cell l47B(g2[45],p2[47],g2[47],p2[45],g3[48],p3[48]);
black_cell l48B(g2[46],p2[48],g2[48],p2[46],g3[49],p3[49]);
black_cell l49B(g2[47],p2[49],g2[49],p2[47],g3[50],p3[50]);
black_cell l50B(g2[48],p2[50],g2[50],p2[48],g3[51],p3[51]);
black_cell l51B(g2[49],p2[51],g2[51],p2[49],g3[52],p3[52]);
black_cell l52B(g2[50],p2[52],g2[52],p2[50],g3[53],p3[53]);
black_cell l53B(g2[51],p2[53],g2[53],p2[51],g3[54],p3[54]);
black_cell l54B(g2[52],p2[54],g2[54],p2[52],g3[55],p3[55]);
black_cell l55B(g2[53],p2[55],g2[55],p2[53],g3[56],p3[56]);
black_cell l56B(g2[54],p2[56],g2[56],p2[54],g3[57],p3[57]);
black_cell l57B(g2[55],p2[57],g2[57],p2[55],g3[58],p3[58]);
black_cell l58B(g2[56],p2[58],g2[58],p2[56],g3[59],p3[59]);
black_cell l59B(g2[57],p2[59],g2[59],p2[57],g3[60],p3[60]);
black_cell l60B(g2[58],p2[60],g2[60],p2[58],g3[61],p3[61]);
black_cell l61B(g2[59],p2[61],g2[61],p2[59],g3[62],p3[62]);
black_cell l62B(g2[60],p2[62],g2[62],p2[60],g3[63],p3[63]);
black_cell l63B(g2[61],p2[63],g2[63],p2[61],g3[64],p3[64]);
//level3
gray_cell l4C(cin[0],p3[4],g3[4],g4[4]);
gray_cell l5C(g2[1],p3[5],g3[5],g4[5]);
gray_cell l6C(g3[2],p3[6],g3[6],g4[6]);
gray_cell l7C(g3[3],p3[7],g3[7],g4[7]);
black_cell l8C(g3[4],p3[8],g3[8],p3[4],g4[8],p4[8]);
black_cell l9C(g3[5],p3[9],g3[9],p3[5],g4[9],p4[9]);
black_cell l10C(g3[6],p3[10],g3[10],p3[6],g4[10],p4[10]);
black_cell l11C(g3[7],p3[11],g3[11],p3[7],g4[11],p4[11]);
black_cell l12C(g3[8],p3[12],g3[12],p3[8],g4[12],p4[12]);
black_cell l13C(g3[9],p3[13],g3[13],p3[9],g4[13],p4[13]);
black_cell l14C(g3[10],p3[14],g3[14],p3[10],g4[14],p4[14]);
black_cell l15C(g3[11],p3[15],g3[15],p3[11],g4[15],p4[15]);
black_cell l16C(g3[12],p3[16],g3[16],p3[12],g4[16],p4[16]);
black_cell l17C(g3[13],p3[17],g3[17],p3[13],g4[17],p4[17]);
black_cell l18C(g3[14],p3[18],g3[18],p3[14],g4[18],p4[18]);
black_cell l19C(g3[15],p3[19],g3[19],p3[15],g4[19],p4[19]);
black_cell l20C(g3[16],p3[20],g3[20],p3[16],g4[20],p4[20]);
black_cell l21C(g3[17],p3[21],g3[21],p3[17],g4[21],p4[21]);
black_cell l22C(g3[18],p3[22],g3[22],p3[18],g4[22],p4[22]);
black_cell l23C(g3[19],p3[23],g3[23],p3[19],g4[23],p4[23]);
black_cell l24C(g3[20],p3[24],g3[24],p3[20],g4[24],p4[24]);
black_cell l25C(g3[21],p3[25],g3[25],p3[21],g4[25],p4[25]);
black_cell l26C(g3[22],p3[26],g3[26],p3[22],g4[26],p4[26]);
black_cell l27C(g3[23],p3[27],g3[27],p3[23],g4[27],p4[27]);
black_cell l28C(g3[24],p3[28],g3[28],p3[24],g4[28],p4[28]);
black_cell l29C(g3[25],p3[29],g3[29],p3[25],g4[29],p4[29]);
black_cell l30C(g3[26],p3[30],g3[30],p3[26],g4[30],p4[30]);
black_cell l31C(g3[27],p3[31],g3[31],p3[27],g4[31],p4[31]);
black_cell l32C(g3[28],p3[32],g3[32],p3[28],g4[32],p4[32]);
black_cell l33C(g3[29],p3[33],g3[33],p3[29],g4[33],p4[33]);
black_cell l34C(g3[30],p3[34],g3[34],p3[30],g4[34],p4[34]);
black_cell l35C(g3[31],p3[35],g3[35],p3[31],g4[35],p4[35]);
black_cell l36C(g3[32],p3[36],g3[36],p3[32],g4[36],p4[36]);
black_cell l37C(g3[33],p3[37],g3[37],p3[33],g4[37],p4[37]);
black_cell l38C(g3[34],p3[38],g3[38],p3[34],g4[38],p4[38]);
black_cell l39C(g3[35],p3[39],g3[39],p3[35],g4[39],p4[39]);
black_cell l40C(g3[36],p3[40],g3[40],p3[36],g4[40],p4[40]);
black_cell l41C(g3[37],p3[41],g3[41],p3[37],g4[41],p4[41]);
black_cell l42C(g3[38],p3[42],g3[42],p3[38],g4[42],p4[42]);
black_cell l43C(g3[39],p3[43],g3[43],p3[39],g4[43],p4[43]);
black_cell l44C(g3[40],p3[44],g3[44],p3[40],g4[44],p4[44]);
black_cell l45C(g3[41],p3[45],g3[45],p3[41],g4[45],p4[45]);
black_cell l46C(g3[42],p3[46],g3[46],p3[42],g4[46],p4[46]);
black_cell l47C(g3[43],p3[47],g3[47],p3[43],g4[47],p4[47]);
black_cell l48C(g3[44],p3[48],g3[48],p3[44],g4[48],p4[48]);
black_cell l49C(g3[45],p3[49],g3[49],p3[45],g4[49],p4[49]);
black_cell l50C(g3[46],p3[50],g3[50],p3[46],g4[50],p4[50]);
black_cell l51C(g3[47],p3[51],g3[51],p3[47],g4[51],p4[51]);
black_cell l52C(g3[48],p3[52],g3[52],p3[48],g4[52],p4[52]);
black_cell l53C(g3[49],p3[53],g3[53],p3[49],g4[53],p4[53]);
black_cell l54C(g3[50],p3[54],g3[54],p3[50],g4[54],p4[54]);
black_cell l55C(g3[51],p3[55],g3[55],p3[51],g4[55],p4[55]);
black_cell l56C(g3[52],p3[56],g3[56],p3[52],g4[56],p4[56]);
black_cell l57C(g3[53],p3[57],g3[57],p3[53],g4[57],p4[57]);
black_cell l58C(g3[54],p3[58],g3[58],p3[54],g4[58],p4[58]);
black_cell l59C(g3[55],p3[59],g3[59],p3[55],g4[59],p4[59]);
black_cell l60C(g3[56],p3[60],g3[60],p3[56],g4[60],p4[60]);
black_cell l61C(g3[57],p3[61],g3[61],p3[57],g4[61],p4[61]);
black_cell l62C(g3[58],p3[62],g3[62],p3[58],g4[62],p4[62]);
black_cell l63C(g3[59],p3[63],g3[63],p3[59],g4[63],p4[63]);
black_cell l64C(g3[60],p3[64],g3[64],p3[60],g4[64],p4[64]);

//level4
gray_cell l8D(cin[0],p4[8],g4[8],g5[8]);
gray_cell l9D(g2[1],p4[9],g4[9],g5[9]);
gray_cell l10D(g3[2],p4[10],g4[10],g5[10]);
gray_cell l11D(g3[3],p4[11],g4[11],g5[11]);
gray_cell l12D(g4[4],p4[12],g4[12],g5[12]);
gray_cell l13D(g4[5],p4[13],g4[13],g5[13]);
gray_cell l14D(g4[6],p4[14],g4[14],g5[14]);
gray_cell l15D(g4[7],p4[15],g4[15],g5[15]);
black_cell l16D(g4[8],p4[16],g4[16],p4[8],g5[16],p5[16]);
black_cell l17D(g4[9],p4[17],g4[17],p4[9],g5[17],p5[17]);
black_cell l18D(g4[10],p4[18],g4[18],p4[10],g5[18],p5[18]);
black_cell l19D(g4[11],p4[19],g4[19],p4[11],g5[19],p5[19]);
black_cell l20D(g4[12],p4[20],g4[20],p4[12],g5[20],p5[20]);
black_cell l21D(g4[13],p4[21],g4[21],p4[13],g5[21],p5[21]);
black_cell l22D(g4[14],p4[22],g4[22],p4[14],g5[22],p5[22]);
black_cell l23D(g4[15],p4[23],g4[23],p4[15],g5[23],p5[23]);
black_cell l24D(g4[16],p4[24],g4[24],p4[16],g5[24],p5[24]);
black_cell l25D(g4[17],p4[25],g4[25],p4[17],g5[25],p5[25]);
black_cell l26D(g4[18],p4[26],g4[26],p4[18],g5[26],p5[26]);
black_cell l27D(g4[19],p4[27],g4[27],p4[19],g5[27],p5[27]);
black_cell l28D(g4[20],p4[28],g4[28],p4[20],g5[28],p5[28]);
black_cell l29D(g4[21],p4[29],g4[29],p4[21],g5[29],p5[29]);
black_cell l30D(g4[22],p4[30],g4[30],p4[22],g5[30],p5[30]);
black_cell l31D(g4[23],p4[31],g4[31],p4[23],g5[31],p5[31]);
black_cell l32D(g4[24],p4[32],g4[32],p4[24],g5[32],p5[32]);
black_cell l33D(g4[25],p4[33],g4[33],p4[25],g5[33],p5[33]);
black_cell l34D(g4[26],p4[34],g4[34],p4[26],g5[34],p5[34]);
black_cell l35D(g4[27],p4[35],g4[35],p4[27],g5[35],p5[35]);
black_cell l36D(g4[28],p4[36],g4[36],p4[28],g5[36],p5[36]);
black_cell l37D(g4[29],p4[37],g4[37],p4[29],g5[37],p5[37]);
black_cell l38D(g4[30],p4[38],g4[38],p4[30],g5[38],p5[38]);
black_cell l39D(g4[31],p4[39],g4[39],p4[31],g5[39],p5[39]);
black_cell l40D(g4[32],p4[40],g4[40],p4[32],g5[40],p5[40]);
black_cell l41D(g4[33],p4[41],g4[41],p4[33],g5[41],p5[41]);
black_cell l42D(g4[34],p4[42],g4[42],p4[34],g5[42],p5[42]);
black_cell l43D(g4[35],p4[43],g4[43],p4[35],g5[43],p5[43]);
black_cell l44D(g4[36],p4[44],g4[44],p4[36],g5[44],p5[44]);
black_cell l45D(g4[37],p4[45],g4[45],p4[37],g5[45],p5[45]);
black_cell l46D(g4[38],p4[46],g4[46],p4[38],g5[46],p5[46]);
black_cell l47D(g4[39],p4[47],g4[47],p4[39],g5[47],p5[47]);
black_cell l48D(g4[40],p4[48],g4[48],p4[40],g5[48],p5[48]);
black_cell l49D(g4[41],p4[49],g4[49],p4[41],g5[49],p5[49]);
black_cell l50D(g4[42],p4[50],g4[50],p4[42],g5[50],p5[50]);
black_cell l51D(g4[43],p4[51],g4[51],p4[43],g5[51],p5[51]);
black_cell l52D(g4[44],p4[52],g4[52],p4[44],g5[52],p5[52]);
black_cell l53D(g4[45],p4[53],g4[53],p4[45],g5[53],p5[53]);
black_cell l54D(g4[46],p4[54],g4[54],p4[46],g5[54],p5[54]);
black_cell l55D(g4[47],p4[55],g4[55],p4[47],g5[55],p5[55]);
black_cell l56D(g4[48],p4[56],g4[56],p4[48],g5[56],p5[56]);
black_cell l57D(g4[49],p4[57],g4[57],p4[49],g5[57],p5[57]);
black_cell l58D(g4[50],p4[58],g4[58],p4[50],g5[58],p5[58]);
black_cell l59D(g4[51],p4[59],g4[59],p4[51],g5[59],p5[59]);
black_cell l60D(g4[52],p4[60],g4[60],p4[52],g5[60],p5[60]);
black_cell l61D(g4[53],p4[61],g4[61],p4[53],g5[61],p5[61]);
black_cell l62D(g4[54],p4[62],g4[62],p4[54],g5[62],p5[62]);
black_cell l63D(g4[55],p4[63],g4[63],p4[55],g5[63],p5[63]);
black_cell l64D(g4[56],p4[64],g4[64],p4[56],g5[64],p5[64]);
//level5
gray_cell l16E(cin[0],p5[16],g5[16],g6[16]);
gray_cell l17E(g2[1],p5[17],g5[17],g6[17]);
gray_cell l18E(g3[2],p5[18],g5[18],g6[18]);
gray_cell l19E(g3[3],p5[19],g5[19],g6[19]);
gray_cell l20E(g4[4],p5[20],g5[20],g6[20]);
gray_cell l21E(g4[5],p5[21],g5[21],g6[21]);
gray_cell l22E(g4[6],p5[22],g5[22],g6[22]);
gray_cell l23E(g4[7],p5[23],g5[23],g6[23]);
gray_cell l24E(g5[8],p5[24],g5[24],g6[24]);
gray_cell l25E(g5[9],p5[25],g5[25],g6[25]);
gray_cell l26E(g5[10],p5[26],g5[26],g6[26]);
gray_cell l27E(g5[11],p5[27],g5[27],g6[27]);
gray_cell l28E(g5[12],p5[28],g5[28],g6[28]);
gray_cell l29E(g5[13],p5[29],g5[29],g6[29]);
gray_cell l30E(g5[14],p5[30],g5[30],g6[30]);
gray_cell l31E(g5[15],p5[31],g5[31],g6[31]);
black_cell l32E(g5[16],p5[32],g5[32],p5[16],g6[32],p6[32]);
black_cell l33E(g5[17],p5[33],g5[33],p5[17],g6[33],p6[33]);
black_cell l34E(g5[18],p5[34],g5[34],p5[18],g6[34],p6[34]);
black_cell l35E(g5[19],p5[35],g5[35],p5[19],g6[35],p6[35]);
black_cell l36E(g5[20],p5[36],g5[36],p5[20],g6[36],p6[36]);
black_cell l37E(g5[21],p5[37],g5[37],p5[21],g6[37],p6[37]);
black_cell l38E(g5[22],p5[38],g5[38],p5[22],g6[38],p6[38]);
black_cell l39E(g5[23],p5[39],g5[39],p5[23],g6[39],p6[39]);
black_cell l40E(g5[24],p5[40],g5[40],p5[24],g6[40],p6[40]);
black_cell l41E(g5[25],p5[41],g5[41],p5[25],g6[41],p6[41]);
black_cell l42E(g5[26],p5[42],g5[42],p5[26],g6[42],p6[42]);
black_cell l43E(g5[27],p5[43],g5[43],p5[27],g6[43],p6[43]);
black_cell l44E(g5[28],p5[44],g5[44],p5[28],g6[44],p6[44]);
black_cell l45E(g5[29],p5[45],g5[45],p5[29],g6[45],p6[45]);
black_cell l46E(g5[30],p5[46],g5[46],p5[30],g6[46],p6[46]);
black_cell l47E(g5[31],p5[47],g5[47],p5[31],g6[47],p6[47]);
black_cell l48E(g5[32],p5[48],g5[48],p5[32],g6[48],p6[48]);
black_cell l49E(g5[33],p5[49],g5[49],p5[33],g6[49],p6[49]);
black_cell l50E(g5[34],p5[50],g5[50],p5[34],g6[50],p6[50]);
black_cell l51E(g5[35],p5[51],g5[51],p5[35],g6[51],p6[51]);
black_cell l52E(g5[36],p5[52],g5[52],p5[36],g6[52],p6[52]);
black_cell l53E(g5[37],p5[53],g5[53],p5[37],g6[53],p6[53]);
black_cell l54E(g5[38],p5[54],g5[54],p5[38],g6[54],p6[54]);
black_cell l55E(g5[39],p5[55],g5[55],p5[39],g6[55],p6[55]);
black_cell l56E(g5[40],p5[56],g5[56],p5[40],g6[56],p6[56]);
black_cell l57E(g5[41],p5[57],g5[57],p5[41],g6[57],p6[57]);
black_cell l58E(g5[42],p5[58],g5[58],p5[42],g6[58],p6[58]);
black_cell l59E(g5[43],p5[59],g5[59],p5[43],g6[59],p6[59]);
black_cell l60E(g5[44],p5[60],g5[60],p5[44],g6[60],p6[60]);
black_cell l61E(g5[45],p5[61],g5[61],p5[45],g6[61],p6[61]);
black_cell l62E(g5[46],p5[62],g5[62],p5[46],g6[62],p6[62]);
black_cell l63E(g5[47],p5[63],g5[63],p5[47],g6[63],p6[63]);
black_cell l64E(g5[48],p5[64],g5[64],p5[48],g6[64],p6[64]);
//LEVEL 6
gray_cell l32F(cin[0],p6[32],g6[32],g7[32]);
gray_cell l33F(g2[1],p6[33],g6[33],g7[33]);
gray_cell l34F(g3[2],p6[34],g6[34],g7[34]);
gray_cell l35F(g3[3],p6[35],g6[35],g7[35]);
gray_cell l36F(g4[4],p6[36],g6[36],g7[36]);
gray_cell l37F(g4[5],p6[37],g6[37],g7[37]);
gray_cell l38F(g4[6],p6[38],g6[38],g7[38]);
gray_cell l39F(g4[7],p6[39],g6[39],g7[39]);
gray_cell l40F(g5[8],p6[40],g6[40],g7[40]);
gray_cell l41F(g5[9],p6[41],g6[41],g7[41]);
gray_cell l42F(g5[10],p6[42],g6[42],g7[42]);
gray_cell l43F(g5[11],p6[43],g6[43],g7[43]);
gray_cell l44F(g5[12],p6[44],g6[44],g7[44]);
gray_cell l45F(g5[13],p6[45],g6[45],g7[45]);
gray_cell l46F(g5[14],p6[46],g6[46],g7[46]);
gray_cell l47F(g5[15],p6[47],g6[47],g7[47]);
gray_cell l48F(g6[16],p6[48],g6[48],g7[48]);
gray_cell l49F(g6[17],p6[59],g6[49],g7[49]);
gray_cell l50F(g6[18],p6[50],g6[50],g7[50]);
gray_cell l51F(g6[19],p6[51],g6[51],g7[51]);
gray_cell l52F(g6[20],p6[52],g6[52],g7[52]);
gray_cell l53F(g6[21],p6[53],g6[53],g7[53]);
gray_cell l54F(g6[22],p6[54],g6[54],g7[54]);
gray_cell l55F(g6[23],p6[55],g6[55],g7[55]);
gray_cell l56F(g6[24],p6[56],g6[56],g7[56]);
gray_cell l57F(g6[25],p6[57],g6[57],g7[57]);
gray_cell l58F(g6[26],p6[58],g6[58],g7[58]);
gray_cell l59F(g6[27],p6[69],g6[59],g7[59]);
gray_cell l60F(g6[28],p6[60],g6[60],g7[60]);
gray_cell l61F(g6[29],p6[61],g6[61],g7[61]);
gray_cell l62F(g6[30],p6[62],g6[62],g7[62]);
gray_cell l63F(g6[31],p6[63],g6[63],g7[63]);
gray_cell l64F(g6[32],p6[64],g6[64],cout);
//xor with and
and_xor lZ0(x[0],y[0],p1[0],g1[0]);
and_xor lZ1(x[1],y[1],p1[1],g1[1]);
and_xor lZ2(x[2],y[2],p1[2],g1[2]);
and_xor lZ3(x[3],y[3],p1[3],g1[3]);
and_xor lZ4(x[4],y[4],p1[4],g1[4]);
and_xor lZ5(x[5],y[5],p1[5],g1[5]);
and_xor lZ6(x[6],y[6],p1[6],g1[6]);
and_xor lZ7(x[7],y[7],p1[7],g1[7]);
and_xor lZ8(x[8],y[8],p1[8],g1[8]);
and_xor lZ9(x[9],y[9],p1[9],g1[9]);
and_xor lZ10(x[10],y[10],p1[10],g1[10]);
and_xor lZ11(x[11],y[11],p1[11],g1[11]);
and_xor lZ12(x[12],y[12],p1[12],g1[12]);
and_xor lZ13(x[13],y[13],p1[13],g1[13]);
and_xor lZ14(x[14],y[14],p1[14],g1[14]);
and_xor lZ15(x[15],y[15],p1[15],g1[15]);
and_xor lZ16(x[16],y[16],p1[16],g1[16]);
and_xor lZ17(x[17],y[17],p1[17],g1[17]);
and_xor lZ18(x[18],y[18],p1[18],g1[18]);
and_xor lZ19(x[19],y[19],p1[19],g1[19]);
and_xor lZ20(x[20],y[20],p1[20],g1[20]);
and_xor lZ21(x[21],y[21],p1[21],g1[21]);
and_xor lZ22(x[22],y[22],p1[22],g1[22]);
and_xor lZ23(x[23],y[23],p1[23],g1[23]);
and_xor lZ24(x[24],y[24],p1[24],g1[24]);
and_xor lZ25(x[25],y[25],p1[25],g1[25]);
and_xor lZ26(x[26],y[26],p1[26],g1[26]);
and_xor lZ27(x[27],y[27],p1[27],g1[27]);
and_xor lZ28(x[28],y[28],p1[28],g1[28]);
and_xor lZ29(x[29],y[29],p1[29],g1[29]);
and_xor lZ30(x[30],y[30],p1[30],g1[30]);
and_xor lZ31(x[31],y[31],p1[31],g1[31]);
and_xor lZ32(x[32],y[32],p1[32],g1[32]);
and_xor lZ33(x[33],y[33],p1[33],g1[33]);
and_xor lZ34(x[34],y[34],p1[34],g1[34]);
and_xor lZ35(x[35],y[35],p1[35],g1[35]);
and_xor lZ36(x[36],y[36],p1[36],g1[36]);
and_xor lZ37(x[37],y[37],p1[37],g1[37]);
and_xor lZ38(x[38],y[38],p1[38],g1[38]);
and_xor lZ39(x[39],y[39],p1[39],g1[39]);
and_xor lZ40(x[40],y[40],p1[40],g1[40]);
and_xor lZ41(x[41],y[41],p1[41],g1[41]);
and_xor lZ42(x[42],y[42],p1[42],g1[42]);
and_xor lZ43(x[43],y[43],p1[43],g1[43]);
and_xor lZ44(x[44],y[44],p1[44],g1[44]);
and_xor lZ45(x[45],y[45],p1[45],g1[45]);
and_xor lZ46(x[46],y[46],p1[46],g1[46]);
and_xor lZ47(x[47],y[47],p1[47],g1[47]);
and_xor lZ48(x[48],y[48],p1[48],g1[48]);
and_xor lZ49(x[49],y[49],p1[49],g1[49]);
and_xor lZ50(x[50],y[50],p1[50],g1[50]);
and_xor lZ51(x[51],y[51],p1[51],g1[51]);
and_xor lZ52(x[52],y[52],p1[52],g1[52]);
and_xor lZ53(x[53],y[53],p1[53],g1[53]);
and_xor lZ54(x[54],y[54],p1[54],g1[54]);
and_xor lZ55(x[55],y[55],p1[55],g1[55]);
and_xor lZ56(x[56],y[56],p1[56],g1[56]);
and_xor lZ57(x[57],y[57],p1[57],g1[57]);
and_xor lZ58(x[58],y[58],p1[58],g1[58]);
and_xor lZ59(x[59],y[59],p1[59],g1[59]);
and_xor lZ60(x[60],y[60],p1[60],g1[60]);
and_xor lZ61(x[61],y[61],p1[61],g1[61]);
and_xor lZ62(x[62],y[62],p1[62],g1[62]);
and_xor lZ63(x[63],y[63],p1[63],g1[63]);

//outputs
xor_1 x1(sum[0],cin[0],p1[0]);
xor_1 x2(sum[1],g2[0],p1[1]);
xor_1 x3(sum[2],g3[2],p1[2]);
xor_1 x4(sum[3],g3[3],p1[3]);
xor_1 x5(sum[4],g4[4],p1[4]);
xor_1 x6(sum[5],g4[5],p1[5]);
xor_1 x7(sum[6],g4[6],p1[6]);
xor_1 x8(sum[7],g4[7],p1[7]);
xor_1 x9(sum[8],g5[8],p1[8]);
xor_1 x10(sum[9],g5[9],p1[9]);
xor_1 x11(sum[10],g5[10],p1[10]);
xor_1 x12(sum[11],g5[11],p1[11]);
xor_1 x13(sum[12],g5[12],p1[12]);
xor_1 x14(sum[13],g5[13],p1[13]);
xor_1 x15(sum[14],g5[14],p1[14]);
xor_1 x16(sum[15],g5[15],p1[15]);
xor_1 x17(sum[16],g6[16],p1[16]);
xor_1 x18(sum[17],g6[17],p1[17]);
xor_1 x19(sum[18],g6[18],p1[18]);
xor_1 x20(sum[19],g6[19],p1[19]);
xor_1 x21(sum[20],g6[20],p1[20]);
xor_1 x22(sum[21],g6[21],p1[21]);
xor_1 x23(sum[22],g6[22],p1[22]);
xor_1 x24(sum[23],g6[23],p1[23]);
xor_1 x25(sum[24],g6[24],p1[24]);
xor_1 x26(sum[25],g6[25],p1[25]);
xor_1 x27(sum[26],g6[26],p1[26]);
xor_1 x28(sum[27],g6[27],p1[27]);
xor_1 x29(sum[28],g6[28],p1[28]);
xor_1 x30(sum[29],g6[29],p1[29]);
xor_1 x31(sum[30],g6[30],p1[30]);
xor_1 x32(sum[31],g6[31],p1[31]);
xor_1 x33(sum[32],g7[32],p1[32]);
xor_1 x34(sum[33],g7[33],p1[33]);
xor_1 x35(sum[34],g7[34],p1[34]);
xor_1 x36(sum[35],g7[35],p1[35]);
xor_1 x37(sum[36],g7[36],p1[36]);
xor_1 x38(sum[37],g7[37],p1[37]);
xor_1 x39(sum[38],g7[38],p1[38]);
xor_1 x40(sum[39],g7[39],p1[39]);
xor_1 x41(sum[40],g7[40],p1[40]);
xor_1 x42(sum[41],g7[41],p1[41]);
xor_1 x43(sum[42],g7[42],p1[42]);
xor_1 x44(sum[43],g7[43],p1[43]);
xor_1 x45(sum[44],g7[44],p1[44]);
xor_1 x46(sum[45],g7[45],p1[45]);
xor_1 x47(sum[46],g7[46],p1[46]);
xor_1 x48(sum[47],g7[47],p1[47]);
xor_1 x49(sum[48],g7[48],p1[48]);
xor_1 x50(sum[49],g7[49],p1[49]);
xor_1 x51(sum[50],g7[50],p1[50]);
xor_1 x52(sum[51],g7[51],p1[51]);
xor_1 x53(sum[52],g7[52],p1[52]);
xor_1 x54(sum[53],g7[53],p1[53]);
xor_1 x55(sum[54],g7[54],p1[54]);
xor_1 x56(sum[55],g7[55],p1[55]);
xor_1 x57(sum[56],g7[56],p1[56]);
xor_1 x58(sum[57],g7[57],p1[57]);
xor_1 x59(sum[58],g7[58],p1[58]);
xor_1 x60(sum[59],g7[59],p1[59]);
xor_1 x61(sum[60],g7[60],p1[60]);
xor_1 x62(sum[61],g7[61],p1[61]);
xor_1 x63(sum[62],g7[62],p1[62]);
xor_1 x64(sum[63],g7[63],p1[63]);
//endmodule declaration
endmodule



//module declaration
module gray_cell(Gkj,Pik,Gik,G);
//port declaration
input Gkj,Pik,Gik;
output G;
wire Y;
//gate instantiation
and(Y,Gkj,Pik);
or(G,Y,Gik);
//endmodule declaration
endmodule



//module declaration
module black_cell(Gkj,Pik,Gik,Pkj,G,P);
//port declaration
input Gkj,Pik,Gik,Pkj;
output G,P;
wire Y;
//gate instantiation
and(Y,Gkj,Pik);
or(G,Gik,Y);
and(P,Pkj,Pik);
//endmodule declaration
endmodule




//module declaration
module and_xor(a,b,p,g);
//port declaration
input a,b;
output p,g;
//gate instantiation
xor(p,a,b);
and(g,a,b);
//endmodule declaration
endmodule


//xor module
module xor_1(y,a,b);
input a,b;
output y;
xor(y,a,b);
endmodule
